module testingModule (
    A,B,X
);

input A; 
input B; 
output X; 

assign X = A & B; 

endmodule